module pro(propegator, a, b);
input a, b;
output propegator;

xor result(propegator, a, b);
endmodule