module gen(generator, a, b);
input a, b;
output generator;
and result(generator, a, b);
endmodule